//top
// `define	  SIM
  `define	  SRC

/*********************************/
`ifdef  SIM
    `define	  VIDEO_320_40
`endif

`ifdef  SRC
    `define	  VIDEO_1280_720
`endif

